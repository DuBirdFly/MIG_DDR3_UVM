typedef uvm_sequencer #(TrAxi) AxiMstrSqrAw;
typedef uvm_sequencer #(TrAxi) AxiMstrSqrW;
typedef uvm_sequencer #(TrAxi) AxiMstrSqrAr;

/*
class AxiMstrSqrAw extends uvm_sequencer #(TrAxi);
    `uvm_component_utils(AxiMstrSqrAw)
    function new(string name = "AxiMstrSqrAw", uvm_component parent);
        super.new(name, parent);
    endfunction
endclass

class AxiMstrSqrW extends uvm_sequencer #(TrAxi);
    `uvm_component_utils(AxiMstrSqrW)
    function new(string name = "AxiMstrSqrW", uvm_component parent);
        super.new(name, parent);
    endfunction
endclass

class AxiMstrSqrAr extends uvm_sequencer #(TrAxi);
    `uvm_component_utils(AxiMstrSqrAr)
    function new(string name = "AxiMstrSqrAr", uvm_component parent);
        super.new(name, parent);
    endfunction
endclass
*/

`ifndef __MEM_CONSTANT_SVH__
    `define __MEM_CONSTANT_SVH__

    `define MEM_DQ_WIDTH        32
    `define MEM_DQS_WIDTH       4
    `define MEM_DM_WIDTH        4

    `define MEM_BA_WIDTH        3
    `define MEM_ROW_WIDTH       13
    `define MEM_COL_WIDTH       10
`endif
